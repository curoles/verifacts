
// comment for module1
module module1;
endmodule
