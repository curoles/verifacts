// define 1
`define MODULE1_SV_DEFINE1 42

// define 2
`define MODULE1_SV_DEFINE2 4242

// comment for module1
module module1;
endmodule
