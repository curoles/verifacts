`define MODULE1_SV_DEFINE1 42

// comment for module1
module module1;
endmodule
